`include "lib/opcodes.v"
`timescale 1ns / 1ps

module ALU
 (input      [`W_OPCODE-1:0]  alu_op,
  input      [`W_CPU-1:0]     A,
  input      [`W_CPU-1:0]     B,
  output reg [`W_CPU-1:0]     R,
  output reg overflow,
  output reg isZero);


  always @* begin
    case(alu_op)
      // math
      `ADD : begin
        {overflow, R} = A + B;
      end
      `ADDU : begin
        {overflow, R} = A + B;
      end
      `SUB : begin
        {overflow, R} = A + ~B;
      end
      `SUBU : begin
        {overflow, R} = A + ~B;
      end
      `SLT : begin
        R = `W_CPU'b0;
        if (A >= B)
        R = `W_CPU'b1;
        overflow = 1'b0;
      end
      `SLTU : begin
        R = `W_CPU'b0;
        if (A >= B)
        R = `W_CPU'b1;
        overflow = 1'b0;
      end
      // shifts
      `SLL : begin
        R = A << B; // TODO make sure this is correct
        overflow = 1'b0;
      end
      `SRL : begin
        R = A >> B;
        overflow = 1'b0;
      end
      `SRA : begin
        R = A >>> B;
        overflow = 1'b0;
      end
      // gates
      `AND : begin
        R = A & B;
        overflow = 1'b0;
      end
      // `NAND : begin
      //   R = ~(A & B);
      //   overflow = 1'b0;
      // end // note: not included in lab4b list or opcodes.v
      `OR : begin
        R = A | B;
        overflow = 1'b0;
      end
      `NOR : begin
        R = ~(A | B);
        overflow = 1'b0;
      end
      `XOR : begin
        R = A ^ B;
        overflow = 1'b0;
      end
      default : begin
        R =  `W_CPU-1'b0; // TODO check this is the right syntax
        overflow = 1'b0;
      end
    endcase
  end
endmodule
